`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:20:03 05/31/2017 
// Design Name: 
// Module Name:    song2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module song2(clk,ifplay,SongData);	
input ifplay;
input clk;
output [4:0]SongData;
reg [9:0]state;
initial state=0;
reg[4:0]YinFu;
assign SongData=YinFu;
always @(posedge clk)
begin
   state = state + 1'b1;	
	if(!ifplay)begin state=0;end
   if(state>576) begin state = 1;end//��ʱ����ʵ��ѭ������
	case(state)
		1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16:YinFu=18;
		17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32:YinFu=15;
		33,34:YinFu=11;
		35:YinFu=13;
		36:YinFu=14;
		37:YinFu=16;
		38:YinFu=14;
		39,40:YinFu=13;
		41,42:YinFu=12;
		43,44:YinFu=13;
		45,46,47,48:YinFu=14;
      49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64:YinFu=21;
		65,66:YinFu=9;
		67,68:YinFu=8;
		69,70:YinFu=9;
		71,72:YinFu=12;
		73,74:YinFu=9;
		75,76:YinFu=8;
		77,78:YinFu=9;
		79,80:YinFu=13;
		81,82:YinFu=9;
		83,84:YinFu=8;
		85,86:YinFu=9;
		87,88:YinFu=14;
		89,90,91,92:YinFu=13;
		93,94,95,96:YinFu=11;
		97,98:YinFu=9;
		99,100:YinFu=8;
		101,102:YinFu=9;
		103,104:YinFu=12;
		105,106:YinFu=9;
		107,108:YinFu=8;
		109,110:YinFu=9;
		111,112:YinFu=13;
		113,114,115,116:YinFu=11;
		117,118,119,120:YinFu=8;
		121,122,123,124,125,126,127,128:YinFu=6;
		
		129,130:YinFu=9;
		131,132:YinFu=8;
		133,134:YinFu=9;
		135,136:YinFu=12;
		137,138:YinFu=9;
		139,140:YinFu=8;
		141,142:YinFu=9;
		143,144:YinFu=13;
		
		145,146:YinFu=9;
		147,148:YinFu=8;
		149,150:YinFu=9;
		151,152:YinFu=14;
		153,154,155,156:YinFu=13;
		157,158,159,160:YinFu=11;
		
		161,162:YinFu=8;
		163,164:YinFu=9;
		165,166,167,168:YinFu=5;
		169,170:YinFu=8;
		171,172:YinFu=9;
		173,174:YinFu=5;
		175,176:YinFu=4;
		
		177,178,179,180:YinFu=5;
		181,182,183,184:YinFu=7;
		185,186,187,188,189,190,191,192:YinFu=4;
		
		193,194:YinFu=5;
		195,196:YinFu=7;
		197,198:YinFu=7;
		199,200:YinFu=8;
		201,202:YinFu=8;
		203,204:YinFu=9;
		205,206:YinFu=9;
		207:YinFu=11;
		208:YinFu=12;
		
		209,210,211,212,213,214:YinFu=11;
		215,216:YinFu=9;
		217,218,219,220,221,222,223,224:YinFu=8;
		
		225,226:YinFu=5;
		227,228:YinFu=7;
		229,230:YinFu=7;
		231,232:YinFu=8;
		233,234:YinFu=8;
		235,236:YinFu=9;
		237,238,239,240:YinFu=9;
		
		241,242,243,244:YinFu=5;
		245,246,247,248,249,250,251,252,253,254,255,256:YinFu=4;
		
		257,258:YinFu=5;
		259,260:YinFu=7;
		261,262:YinFu=7;
		263,264:YinFu=8;
		265,266:YinFu=8;
		267,268:YinFu=9;
		269,270:YinFu=9;
		271:YinFu=11;
		272:YinFu=12;
		
		273,274,275,276,277,278:YinFu=11;
		279,280:YinFu=9;
		281,282,283,284,285,286,287,288:YinFu=8;
		
		289,290:YinFu=8;
		291,292:YinFu=9;
		293,294,295,296:YinFu=5;
		297,298:YinFu=8;
		299,300:YinFu=9;
		301,302:YinFu=5;
		303,304:YinFu=4;
		
		305,306,307,308,309,310,311,312,313,314,315,316:YinFu=5;
		317,318:YinFu=5;
		319,320:YinFu=7;
		
		321,322,323,324,325,326:YinFu=8;
		327,328:YinFu=7;
		329,330,331,332:YinFu=5;
		333,334:YinFu=5;
		335,336:YinFu=7;
		
		337,338,339,340,341,342:YinFu=8;
		343,344:YinFu=7;
		345,346,347,348:YinFu=9;
		349,350:YinFu=9;
		351,352:YinFu=11;
		
		353,354,355,356:YinFu=12;
		357,358:YinFu=12;
		359,360:YinFu=11;
		361,362:YinFu=9;
		363,364:YinFu=8;
		365,366,367,368:YinFu=7;
		
		369,370,371,372:YinFu=8;
		373,374,375,376,377,378,379,380:YinFu=9;
		381,382:YinFu=5;
		383,384:YinFu=7;
		
		385,386,387,388,389,390,391:YinFu=8;
		392:YinFu=7;
		393,394,395,396:YinFu=5;
		397,398:YinFu=5;
		399,400:YinFu=7;
		
		401,402,403,404:YinFu=8;
		405,406,407,408:YinFu=7;
		409:YinFu=8;
		410,411,412,413,414,415,416:YinFu=9;
		
		417,418:YinFu=8;
		419,420:YinFu=9;
		421,422,423,424:YinFu=5;
		425,426:YinFu=8;
		427,428:YinFu=9;
		429,430:YinFu=5;
		431,432:YinFu=4;
		
		433,434,435,436,437,438,439,440,441,442,443,444:YinFu=5;
		445,446:YinFu=9;
		447,448:YinFu=11;
		
		449,450,451,452,453,454:YinFu=14;
		455,456:YinFu=13;
		457,458,459,460:YinFu=9;
		461,462:YinFu=9;
		463,464:YinFu=8;
		
		465,466,467,468:YinFu=7;
		469,470:YinFu=7;
		471,472:YinFu=8;
		473,474,475,476:YinFu=9;
		477,478:YinFu=9;
		479,480:YinFu=8;
		
		481,482,483,484:YinFu=7;
		485,486:YinFu=12;
		487,488:YinFu=14;
		489,490:YinFu=13;
		491,492:YinFu=12;
		493,494:YinFu=11;
		495,496:YinFu=8;
		
		497,498,499,500,501,502,503,504,505,506,507,508:YinFu=9;
		509,510:YinFu=9;
		511,512:YinFu=11;
		
		513,514,515,516,517,518:YinFu=14;
		519,520:YinFu=13;
		521,522,523,524:YinFu=9;
		525,526:YinFu=9;
		527,528:YinFu=8;
		
		529,530,531,532:YinFu=7;
		533,534:YinFu=7;
		535,536:YinFu=8;
		537,538,539,540,541,542,543,544:YinFu=9;
		
		545,546:YinFu=8;
		547,548:YinFu=9;
		549,550,551,552:YinFu=5;
		553,554:YinFu=8;
		555,556:YinFu=9;
		557,558:YinFu=5;
		559,560:YinFu=4;
		
		561,562,563,564,565,566,567,568,569,570,571,572,573,574,575,576:YinFu=5;
	
	default:YinFu=5'b10101;
	endcase
end


endmodule

